--
-- Entity: and2
-- Architecture: structural
-- Author: brianw5
-- Date: 09/17/17
--
library STD;
library IEEE;
use IEEE.std_logic_1164.all;

entity nand2 is

port (
    in1     :   in std_logic;
    in2     :   in std_logic;
    out1    :   out std_logic);
end nand2;

architecture structural of nand2 is

begin

    out1 <= not (in1 and in2);

end structural; 
